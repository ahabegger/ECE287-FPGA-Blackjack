module draw(
input [7:0]seed,
output [7:0]card_code,
output [1:0]suit_code
);

/*
This module will generate a random card 
*/



endmodule
