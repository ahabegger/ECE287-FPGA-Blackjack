module card();











endmodule