module dealer();

endmodule
