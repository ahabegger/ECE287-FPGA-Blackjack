module Blackjack();

endmodule