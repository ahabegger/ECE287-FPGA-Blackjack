module hand(
input [4:0]card_1,
input [4:0]card_2,
output [3:0]value1,
output [3:0]value2
);

always@(*)
begin 
	case(card_code)

	endcase


end

endmodule